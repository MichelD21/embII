library  ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package sorter_pkg is
	type input_type is array (0 to 9) of std_logic_vector(15 downto 0);
end sorter_pkg;